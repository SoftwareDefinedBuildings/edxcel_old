module expmod (
    input [64:0] b,
    input [64:0] e,
    input [64:0] m,
    output [64:0] t
    );

wire input [256:0] b;
wire input [256:0] e;
wire input [256:0] m;
reg output [256:0] t;

integer my_int;

endmodule