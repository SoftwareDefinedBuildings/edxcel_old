module decodeint (
    input clk, 
    input rst,
    input [256:0] s,
    output [256:0] int
    );

wire clk;
wire rst;
wire [256:0] s;
reg [256:0] P;
reg on_curve;

//TODO


endmodule