module slide(
    input clk,
    input rst,
    input valid,
    input [0:32*8-1] a,
    output signed [0:256*8-1] r,
    output done
);


function automatic signed [0:256*8-1] for_body;

input [31:0] i;
input [0:256*8-1] r;

begin: slide_blk
    integer b;
    integer k;
    reg break1;
    reg break2;
    if (r[i*8 +: 8] != 8'sh00) begin
          break1 = 0;
          for (b = 1; b <= 6 && (i + b) < 256; b = b + 1) begin
              if (break1 == 1'b0) begin
                  if (r[(i + b)*8 +: 8] != 8'sd0) begin
                      if (($signed(r[i*8 +: 8]) + $signed(r[(i + b)*8 +: 8] << b)) <= 8'sd15) begin
                          r[i*8 +: 8] = $signed(r[i*8 +: 8]) + $signed(r[(i + b)*8 +: 8] << b);
                          r[(i + b)*8 +: 8] = 8'sd0;
                      end else if ((($signed(r[i*8 +: 8]) - $signed(r[(i + b)*8 +: 8] << b))) >= -8'sd15) begin
                          r[i*8 +: 8] = $signed(r[i*8 +: 8]) - $signed(r[(i + b)*8 +: 8] << b);
                          break2 = 0;
                          for (k = i + b; k < 256; k = k + 1) begin
                              if (break2 == 1'b0) begin
                                  if (r[k*8 +: 8] == 8'sd0) begin
                                      r[k*8 +: 8] = 8'sd1;
                                      break2 = 1;
                                  end
                              end
                              if (break2 == 1'b0) begin
                                  r[k*8 +: 8] = 8'sd0;
                              end
                          end
                      end else begin
                          break1 = 1;
                      end
                  end
              end
          end
      end
      
      for_body = r;
end

endfunction



reg signed [0:256*8-1] rr;
reg rdone;

assign r = rr;
assign done = rdone;

reg [32:0] cycle;
reg [32:0] i;

always @ (posedge clk)
begin
    if (rst == 1'b0) begin
        cycle <= 0;
    end else begin
        rdone <= 0;
        cycle <= cycle + 1;
        
        case (cycle)
            32'd0: begin
                       if (valid == 1'b1)
                       begin
                        rr[0*8 +: 8] <= 8'h01 & (a[(0>>>3)*8 +: 8] >>> (0 & 32'sd7));
                        rr[1*8 +: 8] <= 8'h01 & (a[(1>>>3)*8 +: 8] >>> (1 & 32'sd7));
                        rr[2*8 +: 8] <= 8'h01 & (a[(2>>>3)*8 +: 8] >>> (2 & 32'sd7));
                        rr[3*8 +: 8] <= 8'h01 & (a[(3>>>3)*8 +: 8] >>> (3 & 32'sd7));
                        rr[4*8 +: 8] <= 8'h01 & (a[(4>>>3)*8 +: 8] >>> (4 & 32'sd7));
                        rr[5*8 +: 8] <= 8'h01 & (a[(5>>>3)*8 +: 8] >>> (5 & 32'sd7));
                        rr[6*8 +: 8] <= 8'h01 & (a[(6>>>3)*8 +: 8] >>> (6 & 32'sd7));
                        rr[7*8 +: 8] <= 8'h01 & (a[(7>>>3)*8 +: 8] >>> (7 & 32'sd7));
                        rr[8*8 +: 8] <= 8'h01 & (a[(8>>>3)*8 +: 8] >>> (8 & 32'sd7));
                        rr[9*8 +: 8] <= 8'h01 & (a[(9>>>3)*8 +: 8] >>> (9 & 32'sd7));
                        rr[10*8 +: 8] <= 8'h01 & (a[(10>>>3)*8 +: 8] >>> (10 & 32'sd7));
                        rr[11*8 +: 8] <= 8'h01 & (a[(11>>>3)*8 +: 8] >>> (11 & 32'sd7));
                        rr[12*8 +: 8] <= 8'h01 & (a[(12>>>3)*8 +: 8] >>> (12 & 32'sd7));
                        rr[13*8 +: 8] <= 8'h01 & (a[(13>>>3)*8 +: 8] >>> (13 & 32'sd7));
                        rr[14*8 +: 8] <= 8'h01 & (a[(14>>>3)*8 +: 8] >>> (14 & 32'sd7));
                        rr[15*8 +: 8] <= 8'h01 & (a[(15>>>3)*8 +: 8] >>> (15 & 32'sd7));
                        rr[16*8 +: 8] <= 8'h01 & (a[(16>>>3)*8 +: 8] >>> (16 & 32'sd7));
                        rr[17*8 +: 8] <= 8'h01 & (a[(17>>>3)*8 +: 8] >>> (17 & 32'sd7));
                        rr[18*8 +: 8] <= 8'h01 & (a[(18>>>3)*8 +: 8] >>> (18 & 32'sd7));
                        rr[19*8 +: 8] <= 8'h01 & (a[(19>>>3)*8 +: 8] >>> (19 & 32'sd7));
                        rr[20*8 +: 8] <= 8'h01 & (a[(20>>>3)*8 +: 8] >>> (20 & 32'sd7));
                        rr[21*8 +: 8] <= 8'h01 & (a[(21>>>3)*8 +: 8] >>> (21 & 32'sd7));
                        rr[22*8 +: 8] <= 8'h01 & (a[(22>>>3)*8 +: 8] >>> (22 & 32'sd7));
                        rr[23*8 +: 8] <= 8'h01 & (a[(23>>>3)*8 +: 8] >>> (23 & 32'sd7));
                        rr[24*8 +: 8] <= 8'h01 & (a[(24>>>3)*8 +: 8] >>> (24 & 32'sd7));
                        rr[25*8 +: 8] <= 8'h01 & (a[(25>>>3)*8 +: 8] >>> (25 & 32'sd7));
                        rr[26*8 +: 8] <= 8'h01 & (a[(26>>>3)*8 +: 8] >>> (26 & 32'sd7));
                        rr[27*8 +: 8] <= 8'h01 & (a[(27>>>3)*8 +: 8] >>> (27 & 32'sd7));
                        rr[28*8 +: 8] <= 8'h01 & (a[(28>>>3)*8 +: 8] >>> (28 & 32'sd7));
                        rr[29*8 +: 8] <= 8'h01 & (a[(29>>>3)*8 +: 8] >>> (29 & 32'sd7));
                        rr[30*8 +: 8] <= 8'h01 & (a[(30>>>3)*8 +: 8] >>> (30 & 32'sd7));
                        rr[31*8 +: 8] <= 8'h01 & (a[(31>>>3)*8 +: 8] >>> (31 & 32'sd7));
                        rr[32*8 +: 8] <= 8'h01 & (a[(32>>>3)*8 +: 8] >>> (32 & 32'sd7));
                        rr[33*8 +: 8] <= 8'h01 & (a[(33>>>3)*8 +: 8] >>> (33 & 32'sd7));
                        rr[34*8 +: 8] <= 8'h01 & (a[(34>>>3)*8 +: 8] >>> (34 & 32'sd7));
                        rr[35*8 +: 8] <= 8'h01 & (a[(35>>>3)*8 +: 8] >>> (35 & 32'sd7));
                        rr[36*8 +: 8] <= 8'h01 & (a[(36>>>3)*8 +: 8] >>> (36 & 32'sd7));
                        rr[37*8 +: 8] <= 8'h01 & (a[(37>>>3)*8 +: 8] >>> (37 & 32'sd7));
                        rr[38*8 +: 8] <= 8'h01 & (a[(38>>>3)*8 +: 8] >>> (38 & 32'sd7));
                        rr[39*8 +: 8] <= 8'h01 & (a[(39>>>3)*8 +: 8] >>> (39 & 32'sd7));
                        rr[40*8 +: 8] <= 8'h01 & (a[(40>>>3)*8 +: 8] >>> (40 & 32'sd7));
                        rr[41*8 +: 8] <= 8'h01 & (a[(41>>>3)*8 +: 8] >>> (41 & 32'sd7));
                        rr[42*8 +: 8] <= 8'h01 & (a[(42>>>3)*8 +: 8] >>> (42 & 32'sd7));
                        rr[43*8 +: 8] <= 8'h01 & (a[(43>>>3)*8 +: 8] >>> (43 & 32'sd7));
                        rr[44*8 +: 8] <= 8'h01 & (a[(44>>>3)*8 +: 8] >>> (44 & 32'sd7));
                        rr[45*8 +: 8] <= 8'h01 & (a[(45>>>3)*8 +: 8] >>> (45 & 32'sd7));
                        rr[46*8 +: 8] <= 8'h01 & (a[(46>>>3)*8 +: 8] >>> (46 & 32'sd7));
                        rr[47*8 +: 8] <= 8'h01 & (a[(47>>>3)*8 +: 8] >>> (47 & 32'sd7));
                        rr[48*8 +: 8] <= 8'h01 & (a[(48>>>3)*8 +: 8] >>> (48 & 32'sd7));
                        rr[49*8 +: 8] <= 8'h01 & (a[(49>>>3)*8 +: 8] >>> (49 & 32'sd7));
                        rr[50*8 +: 8] <= 8'h01 & (a[(50>>>3)*8 +: 8] >>> (50 & 32'sd7));
                        rr[51*8 +: 8] <= 8'h01 & (a[(51>>>3)*8 +: 8] >>> (51 & 32'sd7));
                        rr[52*8 +: 8] <= 8'h01 & (a[(52>>>3)*8 +: 8] >>> (52 & 32'sd7));
                        rr[53*8 +: 8] <= 8'h01 & (a[(53>>>3)*8 +: 8] >>> (53 & 32'sd7));
                        rr[54*8 +: 8] <= 8'h01 & (a[(54>>>3)*8 +: 8] >>> (54 & 32'sd7));
                        rr[55*8 +: 8] <= 8'h01 & (a[(55>>>3)*8 +: 8] >>> (55 & 32'sd7));
                        rr[56*8 +: 8] <= 8'h01 & (a[(56>>>3)*8 +: 8] >>> (56 & 32'sd7));
                        rr[57*8 +: 8] <= 8'h01 & (a[(57>>>3)*8 +: 8] >>> (57 & 32'sd7));
                        rr[58*8 +: 8] <= 8'h01 & (a[(58>>>3)*8 +: 8] >>> (58 & 32'sd7));
                        rr[59*8 +: 8] <= 8'h01 & (a[(59>>>3)*8 +: 8] >>> (59 & 32'sd7));
                        rr[60*8 +: 8] <= 8'h01 & (a[(60>>>3)*8 +: 8] >>> (60 & 32'sd7));
                        rr[61*8 +: 8] <= 8'h01 & (a[(61>>>3)*8 +: 8] >>> (61 & 32'sd7));
                        rr[62*8 +: 8] <= 8'h01 & (a[(62>>>3)*8 +: 8] >>> (62 & 32'sd7));
                        rr[63*8 +: 8] <= 8'h01 & (a[(63>>>3)*8 +: 8] >>> (63 & 32'sd7));
                        rr[64*8 +: 8] <= 8'h01 & (a[(64>>>3)*8 +: 8] >>> (64 & 32'sd7));
                        rr[65*8 +: 8] <= 8'h01 & (a[(65>>>3)*8 +: 8] >>> (65 & 32'sd7));
                        rr[66*8 +: 8] <= 8'h01 & (a[(66>>>3)*8 +: 8] >>> (66 & 32'sd7));
                        rr[67*8 +: 8] <= 8'h01 & (a[(67>>>3)*8 +: 8] >>> (67 & 32'sd7));
                        rr[68*8 +: 8] <= 8'h01 & (a[(68>>>3)*8 +: 8] >>> (68 & 32'sd7));
                        rr[69*8 +: 8] <= 8'h01 & (a[(69>>>3)*8 +: 8] >>> (69 & 32'sd7));
                        rr[70*8 +: 8] <= 8'h01 & (a[(70>>>3)*8 +: 8] >>> (70 & 32'sd7));
                        rr[71*8 +: 8] <= 8'h01 & (a[(71>>>3)*8 +: 8] >>> (71 & 32'sd7));
                        rr[72*8 +: 8] <= 8'h01 & (a[(72>>>3)*8 +: 8] >>> (72 & 32'sd7));
                        rr[73*8 +: 8] <= 8'h01 & (a[(73>>>3)*8 +: 8] >>> (73 & 32'sd7));
                        rr[74*8 +: 8] <= 8'h01 & (a[(74>>>3)*8 +: 8] >>> (74 & 32'sd7));
                        rr[75*8 +: 8] <= 8'h01 & (a[(75>>>3)*8 +: 8] >>> (75 & 32'sd7));
                        rr[76*8 +: 8] <= 8'h01 & (a[(76>>>3)*8 +: 8] >>> (76 & 32'sd7));
                        rr[77*8 +: 8] <= 8'h01 & (a[(77>>>3)*8 +: 8] >>> (77 & 32'sd7));
                        rr[78*8 +: 8] <= 8'h01 & (a[(78>>>3)*8 +: 8] >>> (78 & 32'sd7));
                        rr[79*8 +: 8] <= 8'h01 & (a[(79>>>3)*8 +: 8] >>> (79 & 32'sd7));
                        rr[80*8 +: 8] <= 8'h01 & (a[(80>>>3)*8 +: 8] >>> (80 & 32'sd7));
                        rr[81*8 +: 8] <= 8'h01 & (a[(81>>>3)*8 +: 8] >>> (81 & 32'sd7));
                        rr[82*8 +: 8] <= 8'h01 & (a[(82>>>3)*8 +: 8] >>> (82 & 32'sd7));
                        rr[83*8 +: 8] <= 8'h01 & (a[(83>>>3)*8 +: 8] >>> (83 & 32'sd7));
                        rr[84*8 +: 8] <= 8'h01 & (a[(84>>>3)*8 +: 8] >>> (84 & 32'sd7));
                        rr[85*8 +: 8] <= 8'h01 & (a[(85>>>3)*8 +: 8] >>> (85 & 32'sd7));
                        rr[86*8 +: 8] <= 8'h01 & (a[(86>>>3)*8 +: 8] >>> (86 & 32'sd7));
                        rr[87*8 +: 8] <= 8'h01 & (a[(87>>>3)*8 +: 8] >>> (87 & 32'sd7));
                        rr[88*8 +: 8] <= 8'h01 & (a[(88>>>3)*8 +: 8] >>> (88 & 32'sd7));
                        rr[89*8 +: 8] <= 8'h01 & (a[(89>>>3)*8 +: 8] >>> (89 & 32'sd7));
                        rr[90*8 +: 8] <= 8'h01 & (a[(90>>>3)*8 +: 8] >>> (90 & 32'sd7));
                        rr[91*8 +: 8] <= 8'h01 & (a[(91>>>3)*8 +: 8] >>> (91 & 32'sd7));
                        rr[92*8 +: 8] <= 8'h01 & (a[(92>>>3)*8 +: 8] >>> (92 & 32'sd7));
                        rr[93*8 +: 8] <= 8'h01 & (a[(93>>>3)*8 +: 8] >>> (93 & 32'sd7));
                        rr[94*8 +: 8] <= 8'h01 & (a[(94>>>3)*8 +: 8] >>> (94 & 32'sd7));
                        rr[95*8 +: 8] <= 8'h01 & (a[(95>>>3)*8 +: 8] >>> (95 & 32'sd7));
                        rr[96*8 +: 8] <= 8'h01 & (a[(96>>>3)*8 +: 8] >>> (96 & 32'sd7));
                        rr[97*8 +: 8] <= 8'h01 & (a[(97>>>3)*8 +: 8] >>> (97 & 32'sd7));
                        rr[98*8 +: 8] <= 8'h01 & (a[(98>>>3)*8 +: 8] >>> (98 & 32'sd7));
                        rr[99*8 +: 8] <= 8'h01 & (a[(99>>>3)*8 +: 8] >>> (99 & 32'sd7));
                        rr[100*8 +: 8] <= 8'h01 & (a[(100>>>3)*8 +: 8] >>> (100 & 32'sd7));
                        rr[101*8 +: 8] <= 8'h01 & (a[(101>>>3)*8 +: 8] >>> (101 & 32'sd7));
                        rr[102*8 +: 8] <= 8'h01 & (a[(102>>>3)*8 +: 8] >>> (102 & 32'sd7));
                        rr[103*8 +: 8] <= 8'h01 & (a[(103>>>3)*8 +: 8] >>> (103 & 32'sd7));
                        rr[104*8 +: 8] <= 8'h01 & (a[(104>>>3)*8 +: 8] >>> (104 & 32'sd7));
                        rr[105*8 +: 8] <= 8'h01 & (a[(105>>>3)*8 +: 8] >>> (105 & 32'sd7));
                        rr[106*8 +: 8] <= 8'h01 & (a[(106>>>3)*8 +: 8] >>> (106 & 32'sd7));
                        rr[107*8 +: 8] <= 8'h01 & (a[(107>>>3)*8 +: 8] >>> (107 & 32'sd7));
                        rr[108*8 +: 8] <= 8'h01 & (a[(108>>>3)*8 +: 8] >>> (108 & 32'sd7));
                        rr[109*8 +: 8] <= 8'h01 & (a[(109>>>3)*8 +: 8] >>> (109 & 32'sd7));
                        rr[110*8 +: 8] <= 8'h01 & (a[(110>>>3)*8 +: 8] >>> (110 & 32'sd7));
                        rr[111*8 +: 8] <= 8'h01 & (a[(111>>>3)*8 +: 8] >>> (111 & 32'sd7));
                        rr[112*8 +: 8] <= 8'h01 & (a[(112>>>3)*8 +: 8] >>> (112 & 32'sd7));
                        rr[113*8 +: 8] <= 8'h01 & (a[(113>>>3)*8 +: 8] >>> (113 & 32'sd7));
                        rr[114*8 +: 8] <= 8'h01 & (a[(114>>>3)*8 +: 8] >>> (114 & 32'sd7));
                        rr[115*8 +: 8] <= 8'h01 & (a[(115>>>3)*8 +: 8] >>> (115 & 32'sd7));
                        rr[116*8 +: 8] <= 8'h01 & (a[(116>>>3)*8 +: 8] >>> (116 & 32'sd7));
                        rr[117*8 +: 8] <= 8'h01 & (a[(117>>>3)*8 +: 8] >>> (117 & 32'sd7));
                        rr[118*8 +: 8] <= 8'h01 & (a[(118>>>3)*8 +: 8] >>> (118 & 32'sd7));
                        rr[119*8 +: 8] <= 8'h01 & (a[(119>>>3)*8 +: 8] >>> (119 & 32'sd7));
                        rr[120*8 +: 8] <= 8'h01 & (a[(120>>>3)*8 +: 8] >>> (120 & 32'sd7));
                        rr[121*8 +: 8] <= 8'h01 & (a[(121>>>3)*8 +: 8] >>> (121 & 32'sd7));
                        rr[122*8 +: 8] <= 8'h01 & (a[(122>>>3)*8 +: 8] >>> (122 & 32'sd7));
                        rr[123*8 +: 8] <= 8'h01 & (a[(123>>>3)*8 +: 8] >>> (123 & 32'sd7));
                        rr[124*8 +: 8] <= 8'h01 & (a[(124>>>3)*8 +: 8] >>> (124 & 32'sd7));
                        rr[125*8 +: 8] <= 8'h01 & (a[(125>>>3)*8 +: 8] >>> (125 & 32'sd7));
                        rr[126*8 +: 8] <= 8'h01 & (a[(126>>>3)*8 +: 8] >>> (126 & 32'sd7));
                        rr[127*8 +: 8] <= 8'h01 & (a[(127>>>3)*8 +: 8] >>> (127 & 32'sd7));
                        rr[128*8 +: 8] <= 8'h01 & (a[(128>>>3)*8 +: 8] >>> (128 & 32'sd7));
                        rr[129*8 +: 8] <= 8'h01 & (a[(129>>>3)*8 +: 8] >>> (129 & 32'sd7));
                        rr[130*8 +: 8] <= 8'h01 & (a[(130>>>3)*8 +: 8] >>> (130 & 32'sd7));
                        rr[131*8 +: 8] <= 8'h01 & (a[(131>>>3)*8 +: 8] >>> (131 & 32'sd7));
                        rr[132*8 +: 8] <= 8'h01 & (a[(132>>>3)*8 +: 8] >>> (132 & 32'sd7));
                        rr[133*8 +: 8] <= 8'h01 & (a[(133>>>3)*8 +: 8] >>> (133 & 32'sd7));
                        rr[134*8 +: 8] <= 8'h01 & (a[(134>>>3)*8 +: 8] >>> (134 & 32'sd7));
                        rr[135*8 +: 8] <= 8'h01 & (a[(135>>>3)*8 +: 8] >>> (135 & 32'sd7));
                        rr[136*8 +: 8] <= 8'h01 & (a[(136>>>3)*8 +: 8] >>> (136 & 32'sd7));
                        rr[137*8 +: 8] <= 8'h01 & (a[(137>>>3)*8 +: 8] >>> (137 & 32'sd7));
                        rr[138*8 +: 8] <= 8'h01 & (a[(138>>>3)*8 +: 8] >>> (138 & 32'sd7));
                        rr[139*8 +: 8] <= 8'h01 & (a[(139>>>3)*8 +: 8] >>> (139 & 32'sd7));
                        rr[140*8 +: 8] <= 8'h01 & (a[(140>>>3)*8 +: 8] >>> (140 & 32'sd7));
                        rr[141*8 +: 8] <= 8'h01 & (a[(141>>>3)*8 +: 8] >>> (141 & 32'sd7));
                        rr[142*8 +: 8] <= 8'h01 & (a[(142>>>3)*8 +: 8] >>> (142 & 32'sd7));
                        rr[143*8 +: 8] <= 8'h01 & (a[(143>>>3)*8 +: 8] >>> (143 & 32'sd7));
                        rr[144*8 +: 8] <= 8'h01 & (a[(144>>>3)*8 +: 8] >>> (144 & 32'sd7));
                        rr[145*8 +: 8] <= 8'h01 & (a[(145>>>3)*8 +: 8] >>> (145 & 32'sd7));
                        rr[146*8 +: 8] <= 8'h01 & (a[(146>>>3)*8 +: 8] >>> (146 & 32'sd7));
                        rr[147*8 +: 8] <= 8'h01 & (a[(147>>>3)*8 +: 8] >>> (147 & 32'sd7));
                        rr[148*8 +: 8] <= 8'h01 & (a[(148>>>3)*8 +: 8] >>> (148 & 32'sd7));
                        rr[149*8 +: 8] <= 8'h01 & (a[(149>>>3)*8 +: 8] >>> (149 & 32'sd7));
                        rr[150*8 +: 8] <= 8'h01 & (a[(150>>>3)*8 +: 8] >>> (150 & 32'sd7));
                        rr[151*8 +: 8] <= 8'h01 & (a[(151>>>3)*8 +: 8] >>> (151 & 32'sd7));
                        rr[152*8 +: 8] <= 8'h01 & (a[(152>>>3)*8 +: 8] >>> (152 & 32'sd7));
                        rr[153*8 +: 8] <= 8'h01 & (a[(153>>>3)*8 +: 8] >>> (153 & 32'sd7));
                        rr[154*8 +: 8] <= 8'h01 & (a[(154>>>3)*8 +: 8] >>> (154 & 32'sd7));
                        rr[155*8 +: 8] <= 8'h01 & (a[(155>>>3)*8 +: 8] >>> (155 & 32'sd7));
                        rr[156*8 +: 8] <= 8'h01 & (a[(156>>>3)*8 +: 8] >>> (156 & 32'sd7));
                        rr[157*8 +: 8] <= 8'h01 & (a[(157>>>3)*8 +: 8] >>> (157 & 32'sd7));
                        rr[158*8 +: 8] <= 8'h01 & (a[(158>>>3)*8 +: 8] >>> (158 & 32'sd7));
                        rr[159*8 +: 8] <= 8'h01 & (a[(159>>>3)*8 +: 8] >>> (159 & 32'sd7));
                        rr[160*8 +: 8] <= 8'h01 & (a[(160>>>3)*8 +: 8] >>> (160 & 32'sd7));
                        rr[161*8 +: 8] <= 8'h01 & (a[(161>>>3)*8 +: 8] >>> (161 & 32'sd7));
                        rr[162*8 +: 8] <= 8'h01 & (a[(162>>>3)*8 +: 8] >>> (162 & 32'sd7));
                        rr[163*8 +: 8] <= 8'h01 & (a[(163>>>3)*8 +: 8] >>> (163 & 32'sd7));
                        rr[164*8 +: 8] <= 8'h01 & (a[(164>>>3)*8 +: 8] >>> (164 & 32'sd7));
                        rr[165*8 +: 8] <= 8'h01 & (a[(165>>>3)*8 +: 8] >>> (165 & 32'sd7));
                        rr[166*8 +: 8] <= 8'h01 & (a[(166>>>3)*8 +: 8] >>> (166 & 32'sd7));
                        rr[167*8 +: 8] <= 8'h01 & (a[(167>>>3)*8 +: 8] >>> (167 & 32'sd7));
                        rr[168*8 +: 8] <= 8'h01 & (a[(168>>>3)*8 +: 8] >>> (168 & 32'sd7));
                        rr[169*8 +: 8] <= 8'h01 & (a[(169>>>3)*8 +: 8] >>> (169 & 32'sd7));
                        rr[170*8 +: 8] <= 8'h01 & (a[(170>>>3)*8 +: 8] >>> (170 & 32'sd7));
                        rr[171*8 +: 8] <= 8'h01 & (a[(171>>>3)*8 +: 8] >>> (171 & 32'sd7));
                        rr[172*8 +: 8] <= 8'h01 & (a[(172>>>3)*8 +: 8] >>> (172 & 32'sd7));
                        rr[173*8 +: 8] <= 8'h01 & (a[(173>>>3)*8 +: 8] >>> (173 & 32'sd7));
                        rr[174*8 +: 8] <= 8'h01 & (a[(174>>>3)*8 +: 8] >>> (174 & 32'sd7));
                        rr[175*8 +: 8] <= 8'h01 & (a[(175>>>3)*8 +: 8] >>> (175 & 32'sd7));
                        rr[176*8 +: 8] <= 8'h01 & (a[(176>>>3)*8 +: 8] >>> (176 & 32'sd7));
                        rr[177*8 +: 8] <= 8'h01 & (a[(177>>>3)*8 +: 8] >>> (177 & 32'sd7));
                        rr[178*8 +: 8] <= 8'h01 & (a[(178>>>3)*8 +: 8] >>> (178 & 32'sd7));
                        rr[179*8 +: 8] <= 8'h01 & (a[(179>>>3)*8 +: 8] >>> (179 & 32'sd7));
                        rr[180*8 +: 8] <= 8'h01 & (a[(180>>>3)*8 +: 8] >>> (180 & 32'sd7));
                        rr[181*8 +: 8] <= 8'h01 & (a[(181>>>3)*8 +: 8] >>> (181 & 32'sd7));
                        rr[182*8 +: 8] <= 8'h01 & (a[(182>>>3)*8 +: 8] >>> (182 & 32'sd7));
                        rr[183*8 +: 8] <= 8'h01 & (a[(183>>>3)*8 +: 8] >>> (183 & 32'sd7));
                        rr[184*8 +: 8] <= 8'h01 & (a[(184>>>3)*8 +: 8] >>> (184 & 32'sd7));
                        rr[185*8 +: 8] <= 8'h01 & (a[(185>>>3)*8 +: 8] >>> (185 & 32'sd7));
                        rr[186*8 +: 8] <= 8'h01 & (a[(186>>>3)*8 +: 8] >>> (186 & 32'sd7));
                        rr[187*8 +: 8] <= 8'h01 & (a[(187>>>3)*8 +: 8] >>> (187 & 32'sd7));
                        rr[188*8 +: 8] <= 8'h01 & (a[(188>>>3)*8 +: 8] >>> (188 & 32'sd7));
                        rr[189*8 +: 8] <= 8'h01 & (a[(189>>>3)*8 +: 8] >>> (189 & 32'sd7));
                        rr[190*8 +: 8] <= 8'h01 & (a[(190>>>3)*8 +: 8] >>> (190 & 32'sd7));
                        rr[191*8 +: 8] <= 8'h01 & (a[(191>>>3)*8 +: 8] >>> (191 & 32'sd7));
                        rr[192*8 +: 8] <= 8'h01 & (a[(192>>>3)*8 +: 8] >>> (192 & 32'sd7));
                        rr[193*8 +: 8] <= 8'h01 & (a[(193>>>3)*8 +: 8] >>> (193 & 32'sd7));
                        rr[194*8 +: 8] <= 8'h01 & (a[(194>>>3)*8 +: 8] >>> (194 & 32'sd7));
                        rr[195*8 +: 8] <= 8'h01 & (a[(195>>>3)*8 +: 8] >>> (195 & 32'sd7));
                        rr[196*8 +: 8] <= 8'h01 & (a[(196>>>3)*8 +: 8] >>> (196 & 32'sd7));
                        rr[197*8 +: 8] <= 8'h01 & (a[(197>>>3)*8 +: 8] >>> (197 & 32'sd7));
                        rr[198*8 +: 8] <= 8'h01 & (a[(198>>>3)*8 +: 8] >>> (198 & 32'sd7));
                        rr[199*8 +: 8] <= 8'h01 & (a[(199>>>3)*8 +: 8] >>> (199 & 32'sd7));
                        rr[200*8 +: 8] <= 8'h01 & (a[(200>>>3)*8 +: 8] >>> (200 & 32'sd7));
                        rr[201*8 +: 8] <= 8'h01 & (a[(201>>>3)*8 +: 8] >>> (201 & 32'sd7));
                        rr[202*8 +: 8] <= 8'h01 & (a[(202>>>3)*8 +: 8] >>> (202 & 32'sd7));
                        rr[203*8 +: 8] <= 8'h01 & (a[(203>>>3)*8 +: 8] >>> (203 & 32'sd7));
                        rr[204*8 +: 8] <= 8'h01 & (a[(204>>>3)*8 +: 8] >>> (204 & 32'sd7));
                        rr[205*8 +: 8] <= 8'h01 & (a[(205>>>3)*8 +: 8] >>> (205 & 32'sd7));
                        rr[206*8 +: 8] <= 8'h01 & (a[(206>>>3)*8 +: 8] >>> (206 & 32'sd7));
                        rr[207*8 +: 8] <= 8'h01 & (a[(207>>>3)*8 +: 8] >>> (207 & 32'sd7));
                        rr[208*8 +: 8] <= 8'h01 & (a[(208>>>3)*8 +: 8] >>> (208 & 32'sd7));
                        rr[209*8 +: 8] <= 8'h01 & (a[(209>>>3)*8 +: 8] >>> (209 & 32'sd7));
                        rr[210*8 +: 8] <= 8'h01 & (a[(210>>>3)*8 +: 8] >>> (210 & 32'sd7));
                        rr[211*8 +: 8] <= 8'h01 & (a[(211>>>3)*8 +: 8] >>> (211 & 32'sd7));
                        rr[212*8 +: 8] <= 8'h01 & (a[(212>>>3)*8 +: 8] >>> (212 & 32'sd7));
                        rr[213*8 +: 8] <= 8'h01 & (a[(213>>>3)*8 +: 8] >>> (213 & 32'sd7));
                        rr[214*8 +: 8] <= 8'h01 & (a[(214>>>3)*8 +: 8] >>> (214 & 32'sd7));
                        rr[215*8 +: 8] <= 8'h01 & (a[(215>>>3)*8 +: 8] >>> (215 & 32'sd7));
                        rr[216*8 +: 8] <= 8'h01 & (a[(216>>>3)*8 +: 8] >>> (216 & 32'sd7));
                        rr[217*8 +: 8] <= 8'h01 & (a[(217>>>3)*8 +: 8] >>> (217 & 32'sd7));
                        rr[218*8 +: 8] <= 8'h01 & (a[(218>>>3)*8 +: 8] >>> (218 & 32'sd7));
                        rr[219*8 +: 8] <= 8'h01 & (a[(219>>>3)*8 +: 8] >>> (219 & 32'sd7));
                        rr[220*8 +: 8] <= 8'h01 & (a[(220>>>3)*8 +: 8] >>> (220 & 32'sd7));
                        rr[221*8 +: 8] <= 8'h01 & (a[(221>>>3)*8 +: 8] >>> (221 & 32'sd7));
                        rr[222*8 +: 8] <= 8'h01 & (a[(222>>>3)*8 +: 8] >>> (222 & 32'sd7));
                        rr[223*8 +: 8] <= 8'h01 & (a[(223>>>3)*8 +: 8] >>> (223 & 32'sd7));
                        rr[224*8 +: 8] <= 8'h01 & (a[(224>>>3)*8 +: 8] >>> (224 & 32'sd7));
                        rr[225*8 +: 8] <= 8'h01 & (a[(225>>>3)*8 +: 8] >>> (225 & 32'sd7));
                        rr[226*8 +: 8] <= 8'h01 & (a[(226>>>3)*8 +: 8] >>> (226 & 32'sd7));
                        rr[227*8 +: 8] <= 8'h01 & (a[(227>>>3)*8 +: 8] >>> (227 & 32'sd7));
                        rr[228*8 +: 8] <= 8'h01 & (a[(228>>>3)*8 +: 8] >>> (228 & 32'sd7));
                        rr[229*8 +: 8] <= 8'h01 & (a[(229>>>3)*8 +: 8] >>> (229 & 32'sd7));
                        rr[230*8 +: 8] <= 8'h01 & (a[(230>>>3)*8 +: 8] >>> (230 & 32'sd7));
                        rr[231*8 +: 8] <= 8'h01 & (a[(231>>>3)*8 +: 8] >>> (231 & 32'sd7));
                        rr[232*8 +: 8] <= 8'h01 & (a[(232>>>3)*8 +: 8] >>> (232 & 32'sd7));
                        rr[233*8 +: 8] <= 8'h01 & (a[(233>>>3)*8 +: 8] >>> (233 & 32'sd7));
                        rr[234*8 +: 8] <= 8'h01 & (a[(234>>>3)*8 +: 8] >>> (234 & 32'sd7));
                        rr[235*8 +: 8] <= 8'h01 & (a[(235>>>3)*8 +: 8] >>> (235 & 32'sd7));
                        rr[236*8 +: 8] <= 8'h01 & (a[(236>>>3)*8 +: 8] >>> (236 & 32'sd7));
                        rr[237*8 +: 8] <= 8'h01 & (a[(237>>>3)*8 +: 8] >>> (237 & 32'sd7));
                        rr[238*8 +: 8] <= 8'h01 & (a[(238>>>3)*8 +: 8] >>> (238 & 32'sd7));
                        rr[239*8 +: 8] <= 8'h01 & (a[(239>>>3)*8 +: 8] >>> (239 & 32'sd7));
                        rr[240*8 +: 8] <= 8'h01 & (a[(240>>>3)*8 +: 8] >>> (240 & 32'sd7));
                        rr[241*8 +: 8] <= 8'h01 & (a[(241>>>3)*8 +: 8] >>> (241 & 32'sd7));
                        rr[242*8 +: 8] <= 8'h01 & (a[(242>>>3)*8 +: 8] >>> (242 & 32'sd7));
                        rr[243*8 +: 8] <= 8'h01 & (a[(243>>>3)*8 +: 8] >>> (243 & 32'sd7));
                        rr[244*8 +: 8] <= 8'h01 & (a[(244>>>3)*8 +: 8] >>> (244 & 32'sd7));
                        rr[245*8 +: 8] <= 8'h01 & (a[(245>>>3)*8 +: 8] >>> (245 & 32'sd7));
                        rr[246*8 +: 8] <= 8'h01 & (a[(246>>>3)*8 +: 8] >>> (246 & 32'sd7));
                        rr[247*8 +: 8] <= 8'h01 & (a[(247>>>3)*8 +: 8] >>> (247 & 32'sd7));
                        rr[248*8 +: 8] <= 8'h01 & (a[(248>>>3)*8 +: 8] >>> (248 & 32'sd7));
                        rr[249*8 +: 8] <= 8'h01 & (a[(249>>>3)*8 +: 8] >>> (249 & 32'sd7));
                        rr[250*8 +: 8] <= 8'h01 & (a[(250>>>3)*8 +: 8] >>> (250 & 32'sd7));
                        rr[251*8 +: 8] <= 8'h01 & (a[(251>>>3)*8 +: 8] >>> (251 & 32'sd7));
                        rr[252*8 +: 8] <= 8'h01 & (a[(252>>>3)*8 +: 8] >>> (252 & 32'sd7));
                        rr[253*8 +: 8] <= 8'h01 & (a[(253>>>3)*8 +: 8] >>> (253 & 32'sd7));
                        rr[254*8 +: 8] <= 8'h01 & (a[(254>>>3)*8 +: 8] >>> (254 & 32'sd7));
                        rr[255*8 +: 8] <= 8'h01 & (a[(255>>>3)*8 +: 8] >>> (255 & 32'sd7));
                       end
                       else
                       begin
                           cycle <= 0;
                       end
                   end
            32'd1: begin
                        rr <= for_body(0, rr);
                    end
           32'd2: begin
                        rr <= for_body(1, rr);
                    end
           32'd3: begin
                        rr <= for_body(2, rr);
                    end
           32'd4: begin
                        rr <= for_body(3, rr);
                    end
           32'd5: begin
                        rr <= for_body(4, rr);
                    end
           32'd6: begin
                        rr <= for_body(5, rr);
                    end
           32'd7: begin
                        rr <= for_body(6, rr);
                    end
           32'd8: begin
                        rr <= for_body(7, rr);
                    end
           32'd9: begin
                        rr <= for_body(8, rr);
                    end
           32'd10: begin
                        rr <= for_body(9, rr);
                    end
           32'd11: begin
                        rr <= for_body(10, rr);
                    end
           32'd12: begin
                        rr <= for_body(11, rr);
                    end
           32'd13: begin
                        rr <= for_body(12, rr);
                    end
           32'd14: begin
                        rr <= for_body(13, rr);
                    end
           32'd15: begin
                        rr <= for_body(14, rr);
                    end
           32'd16: begin
                        rr <= for_body(15, rr);
                    end
           32'd17: begin
                        rr <= for_body(16, rr);
                    end
           32'd18: begin
                        rr <= for_body(17, rr);
                    end
           32'd19: begin
                        rr <= for_body(18, rr);
                    end
           32'd20: begin
                        rr <= for_body(19, rr);
                    end
           32'd21: begin
                        rr <= for_body(20, rr);
                    end
           32'd22: begin
                        rr <= for_body(21, rr);
                    end
           32'd23: begin
                        rr <= for_body(22, rr);
                    end
           32'd24: begin
                        rr <= for_body(23, rr);
                    end
           32'd25: begin
                        rr <= for_body(24, rr);
                    end
           32'd26: begin
                        rr <= for_body(25, rr);
                    end
           32'd27: begin
                        rr <= for_body(26, rr);
                    end
           32'd28: begin
                        rr <= for_body(27, rr);
                    end
           32'd29: begin
                        rr <= for_body(28, rr);
                    end
           32'd30: begin
                        rr <= for_body(29, rr);
                    end
           32'd31: begin
                        rr <= for_body(30, rr);
                    end
           32'd32: begin
                        rr <= for_body(31, rr);
                    end
           32'd33: begin
                        rr <= for_body(32, rr);
                    end
           32'd34: begin
                        rr <= for_body(33, rr);
                    end
           32'd35: begin
                        rr <= for_body(34, rr);
                    end
           32'd36: begin
                        rr <= for_body(35, rr);
                    end
           32'd37: begin
                        rr <= for_body(36, rr);
                    end
           32'd38: begin
                        rr <= for_body(37, rr);
                    end
           32'd39: begin
                        rr <= for_body(38, rr);
                    end
           32'd40: begin
                        rr <= for_body(39, rr);
                    end
           32'd41: begin
                        rr <= for_body(40, rr);
                    end
           32'd42: begin
                        rr <= for_body(41, rr);
                    end
           32'd43: begin
                        rr <= for_body(42, rr);
                    end
           32'd44: begin
                        rr <= for_body(43, rr);
                    end
           32'd45: begin
                        rr <= for_body(44, rr);
                    end
           32'd46: begin
                        rr <= for_body(45, rr);
                    end
           32'd47: begin
                        rr <= for_body(46, rr);
                    end
           32'd48: begin
                        rr <= for_body(47, rr);
                    end
           32'd49: begin
                        rr <= for_body(48, rr);
                    end
           32'd50: begin
                        rr <= for_body(49, rr);
                    end
           32'd51: begin
                        rr <= for_body(50, rr);
                    end
           32'd52: begin
                        rr <= for_body(51, rr);
                    end
           32'd53: begin
                        rr <= for_body(52, rr);
                    end
           32'd54: begin
                        rr <= for_body(53, rr);
                    end
           32'd55: begin
                        rr <= for_body(54, rr);
                    end
           32'd56: begin
                        rr <= for_body(55, rr);
                    end
           32'd57: begin
                        rr <= for_body(56, rr);
                    end
           32'd58: begin
                        rr <= for_body(57, rr);
                    end
           32'd59: begin
                        rr <= for_body(58, rr);
                    end
           32'd60: begin
                        rr <= for_body(59, rr);
                    end
           32'd61: begin
                        rr <= for_body(60, rr);
                    end
           32'd62: begin
                        rr <= for_body(61, rr);
                    end
           32'd63: begin
                        rr <= for_body(62, rr);
                    end
           32'd64: begin
                        rr <= for_body(63, rr);
                    end
           32'd65: begin
                        rr <= for_body(64, rr);
                    end
           32'd66: begin
                        rr <= for_body(65, rr);
                    end
           32'd67: begin
                        rr <= for_body(66, rr);
                    end
           32'd68: begin
                        rr <= for_body(67, rr);
                    end
           32'd69: begin
                        rr <= for_body(68, rr);
                    end
           32'd70: begin
                        rr <= for_body(69, rr);
                    end
           32'd71: begin
                        rr <= for_body(70, rr);
                    end
           32'd72: begin
                        rr <= for_body(71, rr);
                    end
           32'd73: begin
                        rr <= for_body(72, rr);
                    end
           32'd74: begin
                        rr <= for_body(73, rr);
                    end
           32'd75: begin
                        rr <= for_body(74, rr);
                    end
           32'd76: begin
                        rr <= for_body(75, rr);
                    end
           32'd77: begin
                        rr <= for_body(76, rr);
                    end
           32'd78: begin
                        rr <= for_body(77, rr);
                    end
           32'd79: begin
                        rr <= for_body(78, rr);
                    end
           32'd80: begin
                        rr <= for_body(79, rr);
                    end
           32'd81: begin
                        rr <= for_body(80, rr);
                    end
           32'd82: begin
                        rr <= for_body(81, rr);
                    end
           32'd83: begin
                        rr <= for_body(82, rr);
                    end
           32'd84: begin
                        rr <= for_body(83, rr);
                    end
           32'd85: begin
                        rr <= for_body(84, rr);
                    end
           32'd86: begin
                        rr <= for_body(85, rr);
                    end
           32'd87: begin
                        rr <= for_body(86, rr);
                    end
           32'd88: begin
                        rr <= for_body(87, rr);
                    end
           32'd89: begin
                        rr <= for_body(88, rr);
                    end
           32'd90: begin
                        rr <= for_body(89, rr);
                    end
           32'd91: begin
                        rr <= for_body(90, rr);
                    end
           32'd92: begin
                        rr <= for_body(91, rr);
                    end
           32'd93: begin
                        rr <= for_body(92, rr);
                    end
           32'd94: begin
                        rr <= for_body(93, rr);
                    end
           32'd95: begin
                        rr <= for_body(94, rr);
                    end
           32'd96: begin
                        rr <= for_body(95, rr);
                    end
           32'd97: begin
                        rr <= for_body(96, rr);
                    end
           32'd98: begin
                        rr <= for_body(97, rr);
                    end
           32'd99: begin
                        rr <= for_body(98, rr);
                    end
           32'd100: begin
                        rr <= for_body(99, rr);
                    end
           32'd101: begin
                        rr <= for_body(100, rr);
                    end
           32'd102: begin
                        rr <= for_body(101, rr);
                    end
           32'd103: begin
                        rr <= for_body(102, rr);
                    end
           32'd104: begin
                        rr <= for_body(103, rr);
                    end
           32'd105: begin
                        rr <= for_body(104, rr);
                    end
           32'd106: begin
                        rr <= for_body(105, rr);
                    end
           32'd107: begin
                        rr <= for_body(106, rr);
                    end
           32'd108: begin
                        rr <= for_body(107, rr);
                    end
           32'd109: begin
                        rr <= for_body(108, rr);
                    end
           32'd110: begin
                        rr <= for_body(109, rr);
                    end
           32'd111: begin
                        rr <= for_body(110, rr);
                    end
           32'd112: begin
                        rr <= for_body(111, rr);
                    end
           32'd113: begin
                        rr <= for_body(112, rr);
                    end
           32'd114: begin
                        rr <= for_body(113, rr);
                    end
           32'd115: begin
                        rr <= for_body(114, rr);
                    end
           32'd116: begin
                        rr <= for_body(115, rr);
                    end
           32'd117: begin
                        rr <= for_body(116, rr);
                    end
           32'd118: begin
                        rr <= for_body(117, rr);
                    end
           32'd119: begin
                        rr <= for_body(118, rr);
                    end
           32'd120: begin
                        rr <= for_body(119, rr);
                    end
           32'd121: begin
                        rr <= for_body(120, rr);
                    end
           32'd122: begin
                        rr <= for_body(121, rr);
                    end
           32'd123: begin
                        rr <= for_body(122, rr);
                    end
           32'd124: begin
                        rr <= for_body(123, rr);
                    end
           32'd125: begin
                        rr <= for_body(124, rr);
                    end
           32'd126: begin
                        rr <= for_body(125, rr);
                    end
           32'd127: begin
                        rr <= for_body(126, rr);
                    end
           32'd128: begin
                        rr <= for_body(127, rr);
                    end
           32'd129: begin
                        rr <= for_body(128, rr);
                    end
           32'd130: begin
                        rr <= for_body(129, rr);
                    end
           32'd131: begin
                        rr <= for_body(130, rr);
                    end
           32'd132: begin
                        rr <= for_body(131, rr);
                    end
           32'd133: begin
                        rr <= for_body(132, rr);
                    end
           32'd134: begin
                        rr <= for_body(133, rr);
                    end
           32'd135: begin
                        rr <= for_body(134, rr);
                    end
           32'd136: begin
                        rr <= for_body(135, rr);
                    end
           32'd137: begin
                        rr <= for_body(136, rr);
                    end
           32'd138: begin
                        rr <= for_body(137, rr);
                    end
           32'd139: begin
                        rr <= for_body(138, rr);
                    end
           32'd140: begin
                        rr <= for_body(139, rr);
                    end
           32'd141: begin
                        rr <= for_body(140, rr);
                    end
           32'd142: begin
                        rr <= for_body(141, rr);
                    end
           32'd143: begin
                        rr <= for_body(142, rr);
                    end
           32'd144: begin
                        rr <= for_body(143, rr);
                    end
           32'd145: begin
                        rr <= for_body(144, rr);
                    end
           32'd146: begin
                        rr <= for_body(145, rr);
                    end
           32'd147: begin
                        rr <= for_body(146, rr);
                    end
           32'd148: begin
                        rr <= for_body(147, rr);
                    end
           32'd149: begin
                        rr <= for_body(148, rr);
                    end
           32'd150: begin
                        rr <= for_body(149, rr);
                    end
           32'd151: begin
                        rr <= for_body(150, rr);
                    end
           32'd152: begin
                        rr <= for_body(151, rr);
                    end
           32'd153: begin
                        rr <= for_body(152, rr);
                    end
           32'd154: begin
                        rr <= for_body(153, rr);
                    end
           32'd155: begin
                        rr <= for_body(154, rr);
                    end
           32'd156: begin
                        rr <= for_body(155, rr);
                    end
           32'd157: begin
                        rr <= for_body(156, rr);
                    end
           32'd158: begin
                        rr <= for_body(157, rr);
                    end
           32'd159: begin
                        rr <= for_body(158, rr);
                    end
           32'd160: begin
                        rr <= for_body(159, rr);
                    end
           32'd161: begin
                        rr <= for_body(160, rr);
                    end
           32'd162: begin
                        rr <= for_body(161, rr);
                    end
           32'd163: begin
                        rr <= for_body(162, rr);
                    end
           32'd164: begin
                        rr <= for_body(163, rr);
                    end
           32'd165: begin
                        rr <= for_body(164, rr);
                    end
           32'd166: begin
                        rr <= for_body(165, rr);
                    end
           32'd167: begin
                        rr <= for_body(166, rr);
                    end
           32'd168: begin
                        rr <= for_body(167, rr);
                    end
           32'd169: begin
                        rr <= for_body(168, rr);
                    end
           32'd170: begin
                        rr <= for_body(169, rr);
                    end
           32'd171: begin
                        rr <= for_body(170, rr);
                    end
           32'd172: begin
                        rr <= for_body(171, rr);
                    end
           32'd173: begin
                        rr <= for_body(172, rr);
                    end
           32'd174: begin
                        rr <= for_body(173, rr);
                    end
           32'd175: begin
                        rr <= for_body(174, rr);
                    end
           32'd176: begin
                        rr <= for_body(175, rr);
                    end
           32'd177: begin
                        rr <= for_body(176, rr);
                    end
           32'd178: begin
                        rr <= for_body(177, rr);
                    end
           32'd179: begin
                        rr <= for_body(178, rr);
                    end
           32'd180: begin
                        rr <= for_body(179, rr);
                    end
           32'd181: begin
                        rr <= for_body(180, rr);
                    end
           32'd182: begin
                        rr <= for_body(181, rr);
                    end
           32'd183: begin
                        rr <= for_body(182, rr);
                    end
           32'd184: begin
                        rr <= for_body(183, rr);
                    end
           32'd185: begin
                        rr <= for_body(184, rr);
                    end
           32'd186: begin
                        rr <= for_body(185, rr);
                    end
           32'd187: begin
                        rr <= for_body(186, rr);
                    end
           32'd188: begin
                        rr <= for_body(187, rr);
                    end
           32'd189: begin
                        rr <= for_body(188, rr);
                    end
           32'd190: begin
                        rr <= for_body(189, rr);
                    end
           32'd191: begin
                        rr <= for_body(190, rr);
                    end
           32'd192: begin
                        rr <= for_body(191, rr);
                    end
           32'd193: begin
                        rr <= for_body(192, rr);
                    end
           32'd194: begin
                        rr <= for_body(193, rr);
                    end
           32'd195: begin
                        rr <= for_body(194, rr);
                    end
           32'd196: begin
                        rr <= for_body(195, rr);
                    end
           32'd197: begin
                        rr <= for_body(196, rr);
                    end
           32'd198: begin
                        rr <= for_body(197, rr);
                    end
           32'd199: begin
                        rr <= for_body(198, rr);
                    end
           32'd200: begin
                        rr <= for_body(199, rr);
                    end
           32'd201: begin
                        rr <= for_body(200, rr);
                    end
           32'd202: begin
                        rr <= for_body(201, rr);
                    end
           32'd203: begin
                        rr <= for_body(202, rr);
                    end
           32'd204: begin
                        rr <= for_body(203, rr);
                    end
           32'd205: begin
                        rr <= for_body(204, rr);
                    end
           32'd206: begin
                        rr <= for_body(205, rr);
                    end
           32'd207: begin
                        rr <= for_body(206, rr);
                    end
           32'd208: begin
                        rr <= for_body(207, rr);
                    end
           32'd209: begin
                        rr <= for_body(208, rr);
                    end
           32'd210: begin
                        rr <= for_body(209, rr);
                    end
           32'd211: begin
                        rr <= for_body(210, rr);
                    end
           32'd212: begin
                        rr <= for_body(211, rr);
                    end
           32'd213: begin
                        rr <= for_body(212, rr);
                    end
           32'd214: begin
                        rr <= for_body(213, rr);
                    end
           32'd215: begin
                        rr <= for_body(214, rr);
                    end
           32'd216: begin
                        rr <= for_body(215, rr);
                    end
           32'd217: begin
                        rr <= for_body(216, rr);
                    end
           32'd218: begin
                        rr <= for_body(217, rr);
                    end
           32'd219: begin
                        rr <= for_body(218, rr);
                    end
           32'd220: begin
                        rr <= for_body(219, rr);
                    end
           32'd221: begin
                        rr <= for_body(220, rr);
                    end
           32'd222: begin
                        rr <= for_body(221, rr);
                    end
           32'd223: begin
                        rr <= for_body(222, rr);
                    end
           32'd224: begin
                        rr <= for_body(223, rr);
                    end
           32'd225: begin
                        rr <= for_body(224, rr);
                    end
           32'd226: begin
                        rr <= for_body(225, rr);
                    end
           32'd227: begin
                        rr <= for_body(226, rr);
                    end
           32'd228: begin
                        rr <= for_body(227, rr);
                    end
           32'd229: begin
                        rr <= for_body(228, rr);
                    end
           32'd230: begin
                        rr <= for_body(229, rr);
                    end
           32'd231: begin
                        rr <= for_body(230, rr);
                    end
           32'd232: begin
                        rr <= for_body(231, rr);
                    end
           32'd233: begin
                        rr <= for_body(232, rr);
                    end
           32'd234: begin
                        rr <= for_body(233, rr);
                    end
           32'd235: begin
                        rr <= for_body(234, rr);
                    end
           32'd236: begin
                        rr <= for_body(235, rr);
                    end
           32'd237: begin
                        rr <= for_body(236, rr);
                    end
           32'd238: begin
                        rr <= for_body(237, rr);
                    end
           32'd239: begin
                        rr <= for_body(238, rr);
                    end
           32'd240: begin
                        rr <= for_body(239, rr);
                    end
           32'd241: begin
                        rr <= for_body(240, rr);
                    end
           32'd242: begin
                        rr <= for_body(241, rr);
                    end
           32'd243: begin
                        rr <= for_body(242, rr);
                    end
           32'd244: begin
                        rr <= for_body(243, rr);
                    end
           32'd245: begin
                        rr <= for_body(244, rr);
                    end
           32'd246: begin
                        rr <= for_body(245, rr);
                    end
           32'd247: begin
                        rr <= for_body(246, rr);
                    end
           32'd248: begin
                        rr <= for_body(247, rr);
                    end
           32'd249: begin
                        rr <= for_body(248, rr);
                    end
           32'd250: begin
                        rr <= for_body(249, rr);
                    end
           32'd251: begin
                        rr <= for_body(250, rr);
                    end
           32'd252: begin
                        rr <= for_body(251, rr);
                    end
           32'd253: begin
                        rr <= for_body(252, rr);
                    end
           32'd254: begin
                        rr <= for_body(253, rr);
                    end
           32'd255: begin
                        rr <= for_body(254, rr);
                        rdone <= 1;
                        cycle <= 0;
                    end
        endcase
    end
end
endmodule